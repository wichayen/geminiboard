	library		ieee,std;
	use			ieee.std_logic_1164.all	;
	use			ieee.std_logic_unsigned.all;
	use			ieee.std_logic_arith.all;
	use			ieee.std_logic_misc.all;

--------------------------------------------------------
	
	entity	SYNC_GEN	is
		port	(
				CLK							:	in	std_logic							;
				RST_L						:	in	std_logic							
				
				);
	end	SYNC_GEN;

	architecture	arcSYNC_GEN	of	SYNC_GEN	is
--	------------------------------------------------------------------	--
--	*component															--
--	------------------------------------------------------------------	--
	
--	------------------------------------------------------------------	--
--	*constant	kName						:	size								:=	; -- 
--	------------------------------------------------------------------	--
	
--	------------------------------------------------------------------	--
--	*signal		wName						:	size								:=	; -- 
--	------------------------------------------------------------------	--
	
--====================================================--

--====================================================--
	
--====================================================--

--====================================================--
	begin
	
	process( CLK , RST_L )
	begin
		if ( RST_L = '0' ) then
			
		elsif ( CLK'event and CLK = '1' ) then
			
		end if;
	end process;
	
	
	end	arcSYNC_GEN;
